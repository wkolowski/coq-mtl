(** This module can be used to import/export everything from the directory
    Control/. *)

From CoqMTL Require Export Control.Alternative.
From CoqMTL Require Export Control.Applicative.
From CoqMTL Require Export Control.CommutativeApplicative.
From CoqMTL Require Export Control.Foldable.
From CoqMTL Require Export Control.Functor.
From CoqMTL Require Export Control.Monad.