(** This module exports all monad transformer instances. *)

Require Export Control.Monad.Trans.ContT.
Require Export Control.Monad.Trans.FreeT.
Require Export Control.Monad.Trans.ListT.
Require Export Control.Monad.Trans.OptionT.
Require Export Control.Monad.Trans.ReaderT.
Require Export Control.Monad.Trans.RoseTreeT.
Require Export Control.Monad.Trans.RWST.
Require Export Control.Monad.Trans.StateT.
Require Export Control.Monad.Trans.SumT.
Require Export Control.Monad.Trans.WriterT.