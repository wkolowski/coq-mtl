(** This module exports all monad transformer instances. *)

Require Export HSLib.Control.Monad.Trans.ContT.
Require Export HSLib.Control.Monad.Trans.FreeT.
Require Export HSLib.Control.Monad.Trans.ListT.
Require Export HSLib.Control.Monad.Trans.OptionT.
Require Export HSLib.Control.Monad.Trans.ReaderT.
Require Export HSLib.Control.Monad.Trans.RoseTreeT.
Require Export HSLib.Control.Monad.Trans.RWST.
Require Export HSLib.Control.Monad.Trans.StateT.
Require Export HSLib.Control.Monad.Trans.SumT.
Require Export HSLib.Control.Monad.Trans.WriterT.