(** A module that can be used to important all monadic classes except the
    alternative ones for nondeterminism. *)

Require Export Control.Monad.Class.MonadAlt.
Require Export Control.Monad.Class.MonadExcept.
Require Export Control.Monad.Class.MonadFail.
Require Export Control.Monad.Class.MonadFree.
Require Export Control.Monad.Class.MonadNondet.
Require Export Control.Monad.Class.MonadReader.
Require Export Control.Monad.Class.MonadState.
Require Export Control.Monad.Class.MonadStateNondet.
Require Export Control.Monad.Class.MonadWriter.

(*
Require Export Control.Monad.Class.MonadAlt2.
Require Export Control.Monad.Class.MonadAltSet.
Require Export Control.Monad.Class.MonadAltBag.
*)