(** This module can be used to import/export everything from the directory
    Control/. *)

Require Export Control.Alternative.
Require Export Control.Applicative.
Require Export Control.CommutativeApplicative.
Require Export Control.Foldable.
Require Export Control.Functor.
Require Export Control.Monad.