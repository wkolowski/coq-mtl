(** This module exports all monad transformer instances. *)

From CoqMTL Require Export Control.Monad.Trans.ContT.
From CoqMTL Require Export Control.Monad.Trans.FreeT.
From CoqMTL Require Export Control.Monad.Trans.ListT.
From CoqMTL Require Export Control.Monad.Trans.OptionT.
From CoqMTL Require Export Control.Monad.Trans.ReaderT.
From CoqMTL Require Export Control.Monad.Trans.RoseTreeT.
From CoqMTL Require Export Control.Monad.Trans.RWST.
From CoqMTL Require Export Control.Monad.Trans.StateT.
From CoqMTL Require Export Control.Monad.Trans.SumT.
From CoqMTL Require Export Control.Monad.Trans.WriterT.